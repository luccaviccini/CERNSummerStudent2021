entity T01_HelloWorldTb is
end entity;

architecture sim of T01_HelloWorldTb is
begin

    -- TODO: Create process with Hello World code here

end architecture;