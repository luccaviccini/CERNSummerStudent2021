entity T01_helloworldTB is 
end entity;

architecture sim of T01_helloworldTB is
begin 


	process is 
	begin 
		report "Hello World";
		wait;
	
	end process;


end architecture;

